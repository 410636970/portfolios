`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:45:39 11/27/2019 
// Design Name: 
// Module Name:    Binary2BCD 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Binary2BCD( //13bit
   input [12:0] B,
	output [15:0] P);
	
	wire [68:0] w;
	
	add3 C1(1'b0,B[12],B[11],B[10],w[11],w[2],w[1],w[0]);
	add3 C2(w[2],w[1],w[0],B[9],w[10],w[5],w[4],w[3]);
	add3 C3(w[5],w[4],w[3],B[8],w[9],w[8],w[7],w[6]);
	add3 C4(w[8],w[7],w[6],B[7],w[15],w[14],w[13],w[12]);
	add3 C5(w[14],w[13],w[12],B[6],w[22],w[21],w[20],w[19]);
	
	add3 C6(w[21],w[20],w[19],B[5],w[29],w[28],w[27],w[26]);
	add3 C7(w[28],w[27],w[26],B[4],w[39],w[38],w[37],w[36]);
	add3 C8(w[38],w[37],w[36],B[3],w[50],w[49],w[48],w[47]);
	add3 C9(w[49],w[48],w[47],B[2],w[61],w[60],w[59],w[58]);
	add3 C10(w[60],w[59],w[58],B[1],P[4],P[3],P[2],P[1]);
	
	add3 C11(1'b0,w[11],w[10],w[9],w[35],w[18],w[17],w[16]);
	add3 C12(w[18],w[17],w[16],w[15],w[34],w[25],w[24],w[23]);
	add3 C13(w[25],w[24],w[23],w[22],w[33],w[32],w[31],w[30]);
	add3 C14(w[32],w[31],w[30],w[29],w[43],w[42],w[41],w[40]);
	add3 C15(w[42],w[41],w[40],w[39],w[54],w[53],w[52],w[51]);
	
	add3 C16(w[53],w[52],w[51],w[50],w[65],w[64],w[63],w[62]);
	add3 C17(w[64],w[63],w[62],w[61],P[8],P[7],P[6],P[5]);
	/*add3 C18(1'b0,w[35],w[34],w[33],w[71],w[46],w[45],w[44]);
	add3 C19(w[46],w[45],w[44],w[43],w[70],w[57],w[56],w[55]);
	add3 C20(w[57],w[56],w[55],w[54],w[69],w[68],w[67],w[66]);*/
	add3 C18(1'b0,w[35],w[34],w[33],P[15],w[46],w[45],w[44]);
	add3 C19(w[46],w[45],w[44],w[43],P[14],w[57],w[56],w[55]);
	add3 C20(w[57],w[56],w[55],w[54],P[13],w[68],w[67],w[66]);
	
	add3 C21(w[68],w[67],w[66],w[65],P[12],P[11],P[10],P[9]);
	//add3 C22(1'b0,w[71],w[70],w[69],w[72],P[15],P[14],P[13]);
	
	assign P[0]=B[0];
	
endmodule
